*---------- DMP6023LFG Spice Model ----------
.SUBCKT DMP6023LFG 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.01605 
RS 30 3 0.001 
RG 20 2 4.99 
CGS 2 3 2.839E-009 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 1.75E-009 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 
+ TOX = 6E-008 NSUB = 1E+016 KP = 56.71 KAPPA = 49.86 VTO = -2.33 
.MODEL DCGD D CJO = 8.252E-010 VJ = 1 M = 0.5463 
.MODEL DSUB D IS = 2.343E-010 N = 1.216 RS = 0.003391 BV = 71.9 CJO = 1.513E-010 VJ = 0.1 M = 0.1851 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMP6023LFG Spice Model v1.0 Last Revised 2015/7/7